module hello (
);
    initial begin
        $display ("Hello World");
    end
endmodule